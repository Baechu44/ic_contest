module cross_product (AX, AY, BX, BY, cloclwise);
input	[10:0]	AX, AY, BX, BY;
output			cloclwise;//cloclwise = 1...A cross B 指向裡面
wire	[21:0]	tmp, m1, m2;

multiplier u1 (AX, BY, m1);
multiplier u2 (BX, AY, m2);
assign tmp = m1 - m2;

assign cloclwise = tmp[21];

endmodule


module sub (A, B, S);
input	[19:0]	A, B;
output	[21:0]	S;

wire	[10:0]	S_X, S_Y;

assign S = {S_X, S_Y};

assign S_X = {1'b0, A[19:10]} - {1'b0, B[19:10]};
assign S_Y = {1'b0, A[9:0]}   - {1'b0, B[9:0]};

endmodule

module multiplier(A, B, m);
input  [10:0]  A, B;
output [21:0]  m;
wire   [120:0] T;
wire   [61:0]  U;
wire   [42:0]  W;
wire   [31:1]  X;
wire   [30:1]  Y;
wire           C0;
and a1(T[0], A[0], B[0]);
and a2(T[1], A[1], B[0]);
and a3(T[2], A[2], B[0]);
and a4(T[3], A[3], B[0]);
and a5(T[4], A[4], B[0]);
and a6(T[5], A[5], B[0]);
and a7(T[6], A[6], B[0]);
and a8(T[7], A[7], B[0]);
and a9(T[8], A[8], B[0]);
and a10(T[9], A[9], B[0]);
nand a11(T[10], A[10], B[0]);
and a12(T[11], A[0], B[1]);
and a13(T[12], A[1], B[1]);
and a14(T[13], A[2], B[1]);
and a15(T[14], A[3], B[1]);
and a16(T[15], A[4], B[1]);
and a17(T[16], A[5], B[1]);
and a18(T[17], A[6], B[1]);
and a19(T[18], A[7], B[1]);
and a20(T[19], A[8], B[1]);
and a21(T[20], A[9], B[1]);
nand a22(T[21], A[10], B[1]);
and a23(T[22], A[0], B[2]);
and a24(T[23], A[1], B[2]);
and a25(T[24], A[2], B[2]);
and a26(T[25], A[3], B[2]);
and a27(T[26], A[4], B[2]);
and a28(T[27], A[5], B[2]);
and a29(T[28], A[6], B[2]);
and a30(T[29], A[7], B[2]);
and a31(T[30], A[8], B[2]);
and a32(T[31], A[9], B[2]);
nand a33(T[32], A[10], B[2]);
and a34(T[33], A[0], B[3]);
and a35(T[34], A[1], B[3]);
and a36(T[35], A[2], B[3]);
and a37(T[36], A[3], B[3]);
and a38(T[37], A[4], B[3]);
and a39(T[38], A[5], B[3]);
and a40(T[39], A[6], B[3]);
and a41(T[40], A[7], B[3]);
and a42(T[41], A[8], B[3]);
and a43(T[42], A[9], B[3]);
nand a44(T[43], A[10], B[3]);
and a45(T[44], A[0], B[4]);
and a46(T[45], A[1], B[4]);
and a47(T[46], A[2], B[4]);
and a48(T[47], A[3], B[4]);
and a49(T[48], A[4], B[4]);
and a50(T[49], A[5], B[4]);
and a51(T[50], A[6], B[4]);
and a52(T[51], A[7], B[4]);
and a53(T[52], A[8], B[4]);
and a54(T[53], A[9], B[4]);
nand a55(T[54], A[10], B[4]);
and a56(T[55], A[0], B[5]);
and a57(T[56], A[1], B[5]);
and a58(T[57], A[2], B[5]);
and a59(T[58], A[3], B[5]);
and a60(T[59], A[4], B[5]);
and a61(T[60], A[5], B[5]);
and a62(T[61], A[6], B[5]);
and a63(T[62], A[7], B[5]);
and a64(T[63], A[8], B[5]);
and a65(T[64], A[9], B[5]);
nand a66(T[65], A[10], B[5]);
and a67(T[66], A[0], B[6]);
and a68(T[67], A[1], B[6]);
and a69(T[68], A[2], B[6]);
and a70(T[69], A[3], B[6]);
and a71(T[70], A[4], B[6]);
and a72(T[71], A[5], B[6]);
and a73(T[72], A[6], B[6]);
and a74(T[73], A[7], B[6]);
and a75(T[74], A[8], B[6]);
and a76(T[75], A[9], B[6]);
nand a77(T[76], A[10], B[6]);
and a78(T[77], A[0], B[7]);
and a79(T[78], A[1], B[7]);
and a80(T[79], A[2], B[7]);
and a81(T[80], A[3], B[7]);
and a82(T[81], A[4], B[7]);
and a83(T[82], A[5], B[7]);
and a84(T[83], A[6], B[7]);
and a85(T[84], A[7], B[7]);
and a86(T[85], A[8], B[7]);
and a87(T[86], A[9], B[7]);
nand a88(T[87], A[10], B[7]);
and a89(T[88], A[0], B[8]);
and a90(T[89], A[1], B[8]);
and a91(T[90], A[2], B[8]);
and a92(T[91], A[3], B[8]);
and a93(T[92], A[4], B[8]);
and a94(T[93], A[5], B[8]);
and a95(T[94], A[6], B[8]);
and a96(T[95], A[7], B[8]);
and a97(T[96], A[8], B[8]);
and a98(T[97], A[9], B[8]);
nand a99(T[98], A[10], B[8]);
and a100(T[99], A[0], B[9]);
and a101(T[100], A[1], B[9]);
and a102(T[101], A[2], B[9]);
and a103(T[102], A[3], B[9]);
and a104(T[103], A[4], B[9]);
and a105(T[104], A[5], B[9]);
and a106(T[105], A[6], B[9]);
and a107(T[106], A[7], B[9]);
and a108(T[107], A[8], B[9]);
and a109(T[108], A[9], B[9]);
nand a110(T[109], A[10], B[9]);
nand a111(T[110], A[0], B[10]);
nand a112(T[111], A[1], B[10]);
nand a113(T[112], A[2], B[10]);
nand a114(T[113], A[3], B[10]);
nand a115(T[114], A[4], B[10]);
nand a116(T[115], A[5], B[10]);
nand a117(T[116], A[6], B[10]);
nand a118(T[117], A[7], B[10]);
nand a119(T[118], A[8], B[10]);
nand a120(T[119], A[9], B[10]);
and a121(T[120], A[10], B[10]);
ha ha1(U[0], U[1], T[1], T[11]);//stage0...begin
_233counter counter1(U[3:2], U[4], T[3:2], T[13:12], T[22]);
ha ha2(U[5], U[6], T[23], T[33]);
_233counter counter2(U[8:7], U[9], T[5:4], T[15:14], T[24]);
ha ha3(U[10], U[11], T[34], T[44]);
fa fa1(U[12], U[13], T[25], T[35], T[45]);
_73counter counter3(U[15:14], U[16], T[6], T[16], T[26], T[36], T[46], T[56], T[66]);
_73counter counter4(U[18:17], U[19], T[7], T[17], T[27], T[37], T[47], T[57], T[67]);
_73counter counter5(U[21:20], U[22], T[8], T[18], T[28], T[38], T[48], T[58], T[68]);
ha ha4(U[29], U[30], T[78], T[88]);
_73counter counter6(U[24:23], U[25], T[9], T[19], T[29], T[39], T[49], T[59], T[69]);
_73counter counter7(U[27:26], U[28], T[10], T[20], T[30], T[40], T[50], T[60], T[70]);
_233counter counter8(U[32:31], U[33], T[80:79], T[90:89], T[99]);
ha ha5(U[34], U[35], T[100], T[110]);
_233counter counter9(U[37:36], U[38], T[32:31], T[42:41], T[21]);
_73counter counter10(U[40:39], U[41], T[51], T[61], T[71], T[81], T[91], T[101], T[111]);
_73counter counter11(U[43:42], U[44], T[52], T[62], T[72], T[82], T[92], T[102], T[112]);
_73counter counter12(U[46:45], U[47], T[53], T[63], T[73], T[83], T[93], T[103], T[113]);
_73counter counter13(U[49:48], U[50], T[54], T[64], T[74], T[84], T[94], T[104], T[114]);
_233counter counter14(U[52:51], U[53], T[76:75], T[86:85], T[65]);
_233counter counter15(U[55:54], U[56], T[106:105], T[116:115], T[95]);
_233counter counter16(U[58:57], U[59], T[108:107], T[118:117], T[97]);
ha ha6(U[60], U[61], T[109], T[119]);//stage0...end
ha ha7(W[0], W[1], U[1], U[2]);//stage1...begin
ha ha8(W[2], W[3], U[3], U[5]);
fa fa2(W[4], W[5], U[10], U[7], U[6]);
_233counter counter17(W[7:6], W[8], {U[14], T[55]}, {U[13], U[11]}, U[12]);
_233counter counter18(W[10:9], W[11], {U[18], T[77]}, {U[16], U[17]}, U[15]);
ha ha9(W[12], W[13], U[20], U[29]);
_233counter counter19(W[15:14], W[16], {U[24], U[23]}, {U[22], U[31]}, U[19]);
ha ha10(W[17], W[18], U[30], U[21]);
fa fa3(W[19], W[20], U[34], U[26], U[32]);
_73counter counter20(W[22:21], W[23], 1'b1, U[39], U[36], U[35], U[27], U[33], U[25]);
fa fa4(W[24], W[25], U[37], U[40], U[42]);
_233counter counter21(W[27:26], W[28], {U[48], T[43]}, {U[46], U[45]}, U[38]);
ha ha11(W[29], W[30], U[43], U[41]);
_233counter counter22(W[32:31], W[33], {U[52], U[54]}, {U[50], U[51]}, U[49]);
ha ha12(W[34], W[35], T[96], U[55]);
_233counter counter23(W[37:36], W[38], {T[98], T[87]}, {U[58], U[57]}, U[56]);
ha ha13(W[39], W[40], U[59], U[60]);
ha ha14(W[41], W[42], T[120], U[61]);//stage1...end
ha ha15(X[1], X[2], W[1], W[2]);//stage2...begin
_233counter counter24(X[4:3], X[5], {W[6], U[4]}, {U[8], W[3]}, W[4]);
ha ha16(X[6], X[7], W[7], U[9]);
ha ha17(X[8], X[9], W[8], W[9]);
ha ha18(X[10], X[11], W[10], W[12]);
_233counter counter25(X[13:12], X[14], {W[18], W[17]}, {W[19], W[13]}, W[14]);
_233counter counter26(X[16:15], X[17], {U[28], W[20]}, {W[24], W[16]}, W[21]);
_233counter counter27(X[19:18], X[20], {U[44], W[29]}, {W[30], W[25]}, W[26]);
_233counter counter28(X[22:21], X[23], {W[34], U[47]}, {W[32], W[31]}, W[28]);
fa fa5(X[24], X[25], U[53], W[35], W[36]);
ha ha19(X[26], X[27], W[38], W[39]);
ha ha20(X[28], X[29], W[40], W[41]);
ha ha21(X[30], X[31], W[42], 1'b1);//stage2...end
ha ha22(Y[1], Y[2], X[2], X[3]);//stage3...begin
ha ha23(Y[3], Y[4], X[4], W[5]);
ha ha24(Y[5], Y[6], X[6], X[5]);
ha ha25(Y[7], Y[8], X[7], X[8]);
ha ha26(Y[9], Y[10], X[9], X[10]);
_233counter counter29(Y[12:11], Y[13], {W[15], W[11]}, {X[13], X[11]}, X[12]);
ha ha27(Y[14], Y[15], X[14], X[15]);
ha ha28(Y[16], Y[17], X[16], W[22]);
_233counter counter30(Y[19:18], Y[20], {W[27], W[23]}, {X[19], X[18]}, X[17]);
ha ha29(Y[21], Y[22], X[20], X[21]);
fa fa6(Y[23], Y[24], W[33], X[24], X[23]);
ha ha30(Y[25], Y[26], X[25], W[37]);
ha ha31(Y[27], Y[28], X[27], X[28]);
ha ha32(Y[29], Y[30], X[29], X[30]);//stage3...end
assign m[0]=T[0];//stage4...begin
assign m[1]=U[0];
assign m[2]=W[0];
assign m[3]=X[1];
assign m[4]=Y[1];
ha ha33(m[5], C0, Y[2], Y[3]);
cla16 cla1(m[21:6], , , {Y[28], Y[27], Y[26], Y[24], Y[23], Y[22], Y[20], Y[19], Y[17], Y[15], Y[13], Y[12], Y[10], Y[8], Y[6], Y[4]}, {Y[29], 1'b0, X[26], Y[25], 1'b0, X[22], Y[21], 1'b0, Y[18], Y[16], Y[14], 1'b0, Y[11], Y[9], Y[7], Y[5]}, C0);
endmodule
module ha (Sum, Cout, A, B);
input  A, B;
output Sum, Cout;
wire   Cbar, p;
and a1 (Cout, A, B);
not i1 (Cbar, Cout);
or o1 (p, A, B);
and a2 (Sum, Cbar, p);
endmodule
module fa (Sum, Cout, A, B, Cin);
input  A, B, Cin;
output Sum, Cout;
wire   temp1, g1, g2;
ha ha1 (temp1, g1, A, B);
ha ha2 (Sum, g2, temp1, Cin);
or o1 (Cout, g1, g2);
endmodule
module _233counter (Sum, Cout, A, B, Cin);
input [1:0]  A, B;
input        Cin;
output [1:0] Sum;
output       Cout;
wire         c0;
fa fa1 (Sum[0], c0, A[0], B[0], Cin);
fa fa2 (Sum[1], Cout, A[1], B[1], c0);
endmodule
module _73counter (Sum, Cout, A, B, C, D, E, F, G);
input        A, B, C, D, E, F, G;
output [1:0] Sum;
output       Cout;
wire   [1:0] T0,T1;
fa fa1 (T0[0], T0[1], A, B, C);
fa fa2 (T1[0], T1[1], D, E, F);
_233counter counter (Sum, Cout, T0, T1, G);
endmodule
module cla16 (Sum, G, P, A, B, Cin);
input [15:0]  A, B;
input         Cin;
output [15:0] Sum;
output        G, P;
wire [15:0]   gtemp1, ptemp1, ctemp1;
wire [3:0]    gouta, pouta, ctemp2;
rfa r01 (gtemp1[0], ptemp1[0], Sum[0], A[0], B[0], Cin);
rfa r02 (gtemp1[1], ptemp1[1], Sum[1], A[1], B[1], ctemp1[1]);
rfa r03 (gtemp1[2], ptemp1[2], Sum[2], A[2], B[2], ctemp1[2]);
rfa r04 (gtemp1[3], ptemp1[3], Sum[3], A[3], B[3], ctemp1[3]);
bclg4 b1 (ctemp1[3:0], gouta[0], pouta[0], gtemp1[3:0], ptemp1[3:0], Cin);
rfa r05 (gtemp1[4], ptemp1[4], Sum[4], A[4], B[4], ctemp2[1]);
rfa r06 (gtemp1[5], ptemp1[5], Sum[5], A[5], B[5], ctemp1[5]);
rfa r07 (gtemp1[6], ptemp1[6], Sum[6], A[6], B[6], ctemp1[6]);
rfa r08 (gtemp1[7], ptemp1[7], Sum[7], A[7], B[7], ctemp1[7]);
bclg4 b2 (ctemp1[7:4], gouta[1], pouta[1], gtemp1[7:4], ptemp1[7:4], ctemp2[1]);
rfa r09 (gtemp1[8], ptemp1[8], Sum[8], A[8], B[8], ctemp2[2]);
rfa r10 (gtemp1[9], ptemp1[9], Sum[9], A[9], B[9], ctemp1[9]);
rfa r11 (gtemp1[10], ptemp1[10], Sum[10], A[10], B[10], ctemp1[10]);
rfa r12 (gtemp1[11], ptemp1[11], Sum[11], A[11], B[11], ctemp1[11]);
bclg4 b3 (ctemp1[11:8], gouta[2], pouta[2], gtemp1[11:8], ptemp1[11:8], ctemp2[2]);
rfa r13 (gtemp1[12], ptemp1[12], Sum[12], A[12], B[12], ctemp2[3]);
rfa r14 (gtemp1[13], ptemp1[13], Sum[13], A[13], B[13], ctemp1[13]);
rfa r15 (gtemp1[14], ptemp1[14], Sum[14], A[14], B[14], ctemp1[14]);
rfa r16 (gtemp1[15], ptemp1[15], Sum[15], A[15], B[15], ctemp1[15]);
bclg4 b4 (ctemp1[15:12], gouta[3], pouta[3], gtemp1[15:12], ptemp1[15:12], ctemp2[3]);
bclg4 b5 (ctemp2, G, P, gouta, pouta, Cin);
endmodule
module bclg4 (cout, gout, pout, g, p, cin);
input [3:0]  g, p;
input        cin;
output [3:0] cout;
output       gout, pout;
wire         s1, s2, s3, s4, s5, s6, t1, t2, t3;
and a1 (s1, p[0], cin);
or o1 (cout[1], g[0], s1);
and a2 (s2, p[1], g[0]);
and a3 (s3, p[1], p[0], cin);
or o2 (cout[2], g[1], s2, s3);
and a4 (s4, p[2], g[1]);
and a5 (s5, p[2], p[1], g[0]);
and a6 (s6, p[2], p[1], p[0], cin);
or o3 (cout[3], g[2], s4, s5, s6);
and a7 (t1, p[3], g[2]);
and a8 (t2, p[3], p[2], g[1]);
and a9 (t3, p[3], p[2], p[1], g[0]);
or o4 (gout, g[3], t1, t2, t3);
and a10 (pout, p[3], p[2], p[1], p[0]);
endmodule
module rfa (g, p, Sum, A, B, Cin);
input  A, B, Cin;
output Sum, g, p;
wire   s1, gbar;
and a1 (g, A, B);
not i1 (gbar, g);
or o1 (p, A, B);
and a2 (s1, gbar, p);
ha ha1 (Sum, , s1, Cin);
endmodule
